module and1(input b0,b1, output s0);
	assign s0 = b0 & b1;
endmodule